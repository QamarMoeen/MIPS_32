library verilog;
use verilog.vl_types.all;
entity execute_vlg_vec_tst is
end execute_vlg_vec_tst;
