library verilog;
use verilog.vl_types.all;
entity wrapper_vlg_vec_tst is
end wrapper_vlg_vec_tst;
